-------------------------------------------------------------------------------
--
-- Title       : bin_to_ascii
-- Design      : bin_to_ascii
-- Author      : josuesov115@outlook.es
-- Company     : josjos115
--
-------------------------------------------------------------------------------
--
-- File        : bin_to_ascii.vhd
-- Generated   : Mon Dec  7 14:12:11 2020
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.20
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {bin_to_ascii} architecture {bin_to_ascii}}

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity bin_to_ascii is
	port(din : in std_logic_vector(8 downto 0);
	signo : out std_logic_vector(7 downto 0);
	decena : out std_logic_vector(7 downto 0);
	unidad : out std_logic_vector(7 downto 0);
	decima : out std_logic_vector(7 downto 0);
	centesima : out std_logic_vector(7 downto 0));
end bin_to_ascii;

--}} End of automatically maintained section

architecture synth  of bin_to_ascii is
begin
	 with din(8) select signo <=
	"00101011" when '0',			-- signo +
	"00101101" when others;			-- signo -
	
	with din(7 downto 2) select decena <=
	"00110000" when "000000",	--inicia 0
	"00110000" when "000001",
	"00110000" when "000010",
	"00110000" when "000011",
	"00110000" when "000100",
	"00110000" when "000101",
	"00110000" when "000110",
	"00110000" when "000111",
	"00110000" when "001000",
	"00110000" when "001001",
	"00110001" when "001010",	--inicia 1
	"00110001" when "001011",
	"00110001" when "001100",
	"00110001" when "001101",
	"00110001" when "001110",
	"00110001" when "001111",
	"00110001" when "010000",
	"00110001" when "010001",
	"00110001" when "010010",
	"00110001" when "010011",
	"00110010" when "010100",	--inicia 2
	"00110010" when "010101",
	"00110010" when "010110",
	"00110010" when "010111",
	"00110010" when "011000",
	"00110010" when "011001",
	"00110010" when "011010",
	"00110010" when "011011",
	"00110010" when "011100",
	"00110010" when "011101",
	"00110011" when "011110",	--inicia 3
	"00110011" when "011111",
	"00110011" when "100000",	
	"00110011" when "100001",
	"00110011" when "100010",
	"00110011" when "100011",
	"00110011" when "100100",
	"00110011" when "100101",
	"00110011" when "100110",
	"00110011" when "100111",
	"00110100" when "101000",	--inicia 4
	"00110100" when "101001",
	"00110100" when "101010",	
	"00110100" when "101011",
	"00110100" when "101100",
	"00110100" when "101101",
	"00110100" when "101110",
	"00110100" when "101111",
	"00110100" when "110000",
	"00110100" when "110001",
	"00110101" when "110010",	--inicia 5
	"00110101" when "110011",
	"00110101" when "110100",	
	"00110101" when "110101",
	"00110101" when "110110",
	"00110101" when "110111",
	"00110101" when "111000",
	"00110101" when "111001",
	"00110101" when "111010",
	"00110101" when "111011",
	"00110110" when "111100",	--inicia 6
	"00110110" when "111101",
	"00110110" when "111110",	
	"00110110" when others;
	
	
	with din(7 downto 2) select unidad <=
	"00110000" when "000000",	--0
	"00110001" when "000001",	--1
	"00110010" when "000010",	--2
	"00110011" when "000011",	--3
	"00110100" when "000100",    --4
	"00110101" when "000101",    --5
	"00110110" when "000110",    --6
	"00110111" when "000111",    --7
	"00111000" when "001000",    --8
	"00111001" when "001001",    --9
	"00110000" when "001010",    --0
	"00110001" when "001011",    --1
	"00110010" when "001100",    --2
	"00110011" when "001101",    --3
	"00110100" when "001110",    --4
	"00110101" when "001111",    --5
	"00110110" when "010000",    --6
	"00110111" when "010001",    --7
	"00111000" when "010010",    --8
	"00111001" when "010011",    --9
	"00110000" when "010100",    --0
	"00110001" when "010101",
	"00110010" when "010110",
	"00110011" when "010111",
	"00110100" when "011000",
	"00110101" when "011001",
	"00110110" when "011010",
	"00110111" when "011011",
	"00111000" when "011100",
	"00111001" when "011101",
	"00110000" when "011110",
	"00110001" when "011111",
	"00110010" when "100000",	--2
	"00110011" when "100001",	--3
	"00110100" when "100010",	--4
	"00110101" when "100011",	--5
	"00110110" when "100100",    --6
	"00110111" when "100101",    --7
	"00111000" when "100110",    --8
	"00111001" when "100111",    --9
	"00110000" when "101000",    --0
	"00110001" when "101001",    --1
	"00110010" when "101010",    --2
	"00110011" when "101011",    --3
	"00110100" when "101100",    --4
	"00110101" when "101101",    --5
	"00110110" when "101110",    --6
	"00110111" when "101111",    --7
	"00111000" when "110000",    --8
	"00111001" when "110001",    --9
	"00110000" when "110010",    --0
	"00110001" when "110011",    --1
	"00110010" when "110100",    --2
	"00110011" when "110101",
	"00110100" when "110110",
	"00110101" when "110111",
	"00110110" when "111000",
	"00110111" when "111001",
	"00111000" when "111010",
	"00111001" when "111011",
	"00110000" when "111100",
	"00110001" when "111101",
	"00110010" when "111110",
	"00110011" when others;
	
	with din(1 downto 0) select decima <=
	"00110000" when "00",
	"00110010" when "01",
	"00110101" when "10",
	"00110111" when others;
	
	with din(1 downto 0) select centesima <=
	"00110000" when "00",
	"00110101" when "01",
	"00110000" when "10",
	"00110101" when others;
	
end synth;